// Module 